
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h111ef008;
    ram_cell[       1] = 32'h0;  // 32'h5062b5a8;
    ram_cell[       2] = 32'h0;  // 32'hf234ad08;
    ram_cell[       3] = 32'h0;  // 32'h89257f33;
    ram_cell[       4] = 32'h0;  // 32'hb66a0cdf;
    ram_cell[       5] = 32'h0;  // 32'h2fdc72fc;
    ram_cell[       6] = 32'h0;  // 32'h30eca41b;
    ram_cell[       7] = 32'h0;  // 32'hb1c120de;
    ram_cell[       8] = 32'h0;  // 32'hf625243f;
    ram_cell[       9] = 32'h0;  // 32'h5b4d3964;
    ram_cell[      10] = 32'h0;  // 32'h3d8d34a9;
    ram_cell[      11] = 32'h0;  // 32'h30718281;
    ram_cell[      12] = 32'h0;  // 32'h401c03dd;
    ram_cell[      13] = 32'h0;  // 32'h5760629e;
    ram_cell[      14] = 32'h0;  // 32'hed0dd6b2;
    ram_cell[      15] = 32'h0;  // 32'h79c00ca3;
    ram_cell[      16] = 32'h0;  // 32'h8e4a7d97;
    ram_cell[      17] = 32'h0;  // 32'hcda66b04;
    ram_cell[      18] = 32'h0;  // 32'h6cadf6b4;
    ram_cell[      19] = 32'h0;  // 32'h8c240dac;
    ram_cell[      20] = 32'h0;  // 32'hfdd07b19;
    ram_cell[      21] = 32'h0;  // 32'h873598e9;
    ram_cell[      22] = 32'h0;  // 32'h3c2dd510;
    ram_cell[      23] = 32'h0;  // 32'h3d16609f;
    ram_cell[      24] = 32'h0;  // 32'h7073b9f7;
    ram_cell[      25] = 32'h0;  // 32'h662b04bf;
    ram_cell[      26] = 32'h0;  // 32'h3f7b0ab6;
    ram_cell[      27] = 32'h0;  // 32'h99ecef21;
    ram_cell[      28] = 32'h0;  // 32'hf9296db2;
    ram_cell[      29] = 32'h0;  // 32'h91156933;
    ram_cell[      30] = 32'h0;  // 32'h23870f87;
    ram_cell[      31] = 32'h0;  // 32'h395ebba6;
    ram_cell[      32] = 32'h0;  // 32'hec913769;
    ram_cell[      33] = 32'h0;  // 32'ha0e32a17;
    ram_cell[      34] = 32'h0;  // 32'h4e68aa20;
    ram_cell[      35] = 32'h0;  // 32'h8afbfec5;
    ram_cell[      36] = 32'h0;  // 32'h357eafff;
    ram_cell[      37] = 32'h0;  // 32'h2f1ea264;
    ram_cell[      38] = 32'h0;  // 32'he852ffb6;
    ram_cell[      39] = 32'h0;  // 32'hf2ef565d;
    ram_cell[      40] = 32'h0;  // 32'hebc7f75e;
    ram_cell[      41] = 32'h0;  // 32'h3a872ce1;
    ram_cell[      42] = 32'h0;  // 32'hfc75c69d;
    ram_cell[      43] = 32'h0;  // 32'h0c7b6d29;
    ram_cell[      44] = 32'h0;  // 32'ha28c52fb;
    ram_cell[      45] = 32'h0;  // 32'h8d1a5632;
    ram_cell[      46] = 32'h0;  // 32'h0cf68f74;
    ram_cell[      47] = 32'h0;  // 32'h01db3b59;
    ram_cell[      48] = 32'h0;  // 32'h6a2ffc96;
    ram_cell[      49] = 32'h0;  // 32'hb43fdf0a;
    ram_cell[      50] = 32'h0;  // 32'h6901a6ab;
    ram_cell[      51] = 32'h0;  // 32'h9c1425c5;
    ram_cell[      52] = 32'h0;  // 32'hfaed6478;
    ram_cell[      53] = 32'h0;  // 32'hc1b0a6b4;
    ram_cell[      54] = 32'h0;  // 32'ha1ec0c6b;
    ram_cell[      55] = 32'h0;  // 32'he66609f2;
    ram_cell[      56] = 32'h0;  // 32'h3da2d0d5;
    ram_cell[      57] = 32'h0;  // 32'h15c9e7cc;
    ram_cell[      58] = 32'h0;  // 32'hfbdb7d6e;
    ram_cell[      59] = 32'h0;  // 32'h631f0f77;
    ram_cell[      60] = 32'h0;  // 32'h68d4b555;
    ram_cell[      61] = 32'h0;  // 32'h5f3056fd;
    ram_cell[      62] = 32'h0;  // 32'hb5d84a2a;
    ram_cell[      63] = 32'h0;  // 32'h26908903;
    ram_cell[      64] = 32'h0;  // 32'hf65cec55;
    ram_cell[      65] = 32'h0;  // 32'hbed7f028;
    ram_cell[      66] = 32'h0;  // 32'h53761cb1;
    ram_cell[      67] = 32'h0;  // 32'hf7e28506;
    ram_cell[      68] = 32'h0;  // 32'h775ebc52;
    ram_cell[      69] = 32'h0;  // 32'hc74e3fd2;
    ram_cell[      70] = 32'h0;  // 32'hacf67c2c;
    ram_cell[      71] = 32'h0;  // 32'h070e8fed;
    ram_cell[      72] = 32'h0;  // 32'h25a64bab;
    ram_cell[      73] = 32'h0;  // 32'h35b89a81;
    ram_cell[      74] = 32'h0;  // 32'h2ce2f34e;
    ram_cell[      75] = 32'h0;  // 32'h92a53465;
    ram_cell[      76] = 32'h0;  // 32'haa46a213;
    ram_cell[      77] = 32'h0;  // 32'h23561f9d;
    ram_cell[      78] = 32'h0;  // 32'h0d37b6a8;
    ram_cell[      79] = 32'h0;  // 32'ha0f7510f;
    ram_cell[      80] = 32'h0;  // 32'hec9af09a;
    ram_cell[      81] = 32'h0;  // 32'h68a7c715;
    ram_cell[      82] = 32'h0;  // 32'h02e3a596;
    ram_cell[      83] = 32'h0;  // 32'hc15ee4be;
    ram_cell[      84] = 32'h0;  // 32'he6f45fb3;
    ram_cell[      85] = 32'h0;  // 32'h1fb8c2a7;
    ram_cell[      86] = 32'h0;  // 32'h353086a0;
    ram_cell[      87] = 32'h0;  // 32'h8c773ecd;
    ram_cell[      88] = 32'h0;  // 32'he8b24c65;
    ram_cell[      89] = 32'h0;  // 32'hbaf32d7e;
    ram_cell[      90] = 32'h0;  // 32'h5e397e0e;
    ram_cell[      91] = 32'h0;  // 32'h980db751;
    ram_cell[      92] = 32'h0;  // 32'h6f34a226;
    ram_cell[      93] = 32'h0;  // 32'h1adff5eb;
    ram_cell[      94] = 32'h0;  // 32'hdc251a18;
    ram_cell[      95] = 32'h0;  // 32'h17ccf163;
    ram_cell[      96] = 32'h0;  // 32'hc13b8a7e;
    ram_cell[      97] = 32'h0;  // 32'h51bf3fec;
    ram_cell[      98] = 32'h0;  // 32'h62d174b5;
    ram_cell[      99] = 32'h0;  // 32'h4c13be77;
    ram_cell[     100] = 32'h0;  // 32'h12008efd;
    ram_cell[     101] = 32'h0;  // 32'h68a2b6ba;
    ram_cell[     102] = 32'h0;  // 32'haa003ff2;
    ram_cell[     103] = 32'h0;  // 32'hf51e44ad;
    ram_cell[     104] = 32'h0;  // 32'h654921af;
    ram_cell[     105] = 32'h0;  // 32'h750c7a03;
    ram_cell[     106] = 32'h0;  // 32'h692b96d6;
    ram_cell[     107] = 32'h0;  // 32'h97d3343c;
    ram_cell[     108] = 32'h0;  // 32'hd2897f09;
    ram_cell[     109] = 32'h0;  // 32'hd6fba2fc;
    ram_cell[     110] = 32'h0;  // 32'hd4acabe0;
    ram_cell[     111] = 32'h0;  // 32'hd01b81e5;
    ram_cell[     112] = 32'h0;  // 32'hd3d206fb;
    ram_cell[     113] = 32'h0;  // 32'h51965dd6;
    ram_cell[     114] = 32'h0;  // 32'h31af4e89;
    ram_cell[     115] = 32'h0;  // 32'h7584ddb4;
    ram_cell[     116] = 32'h0;  // 32'hcba88545;
    ram_cell[     117] = 32'h0;  // 32'h5643269d;
    ram_cell[     118] = 32'h0;  // 32'he37c9d74;
    ram_cell[     119] = 32'h0;  // 32'h93a0a7ab;
    ram_cell[     120] = 32'h0;  // 32'h22fd9500;
    ram_cell[     121] = 32'h0;  // 32'h9d31c64b;
    ram_cell[     122] = 32'h0;  // 32'h81ca03d2;
    ram_cell[     123] = 32'h0;  // 32'h1d787c4d;
    ram_cell[     124] = 32'h0;  // 32'hacff6980;
    ram_cell[     125] = 32'h0;  // 32'h0c918984;
    ram_cell[     126] = 32'h0;  // 32'h5c842ec8;
    ram_cell[     127] = 32'h0;  // 32'h67c77069;
    ram_cell[     128] = 32'h0;  // 32'h6461f193;
    ram_cell[     129] = 32'h0;  // 32'h3f368823;
    ram_cell[     130] = 32'h0;  // 32'h7808a5a4;
    ram_cell[     131] = 32'h0;  // 32'h3d752c52;
    ram_cell[     132] = 32'h0;  // 32'hd57778a0;
    ram_cell[     133] = 32'h0;  // 32'h173108f4;
    ram_cell[     134] = 32'h0;  // 32'hbcbebb8f;
    ram_cell[     135] = 32'h0;  // 32'hbf49b2af;
    ram_cell[     136] = 32'h0;  // 32'h1e3fb6e2;
    ram_cell[     137] = 32'h0;  // 32'h235c1718;
    ram_cell[     138] = 32'h0;  // 32'hdfb02c9b;
    ram_cell[     139] = 32'h0;  // 32'h0a7e4df3;
    ram_cell[     140] = 32'h0;  // 32'hca166419;
    ram_cell[     141] = 32'h0;  // 32'hefbeb3bd;
    ram_cell[     142] = 32'h0;  // 32'h2f1ade83;
    ram_cell[     143] = 32'h0;  // 32'h12989b9e;
    ram_cell[     144] = 32'h0;  // 32'h828d09b8;
    ram_cell[     145] = 32'h0;  // 32'h456883ba;
    ram_cell[     146] = 32'h0;  // 32'ha6597965;
    ram_cell[     147] = 32'h0;  // 32'h2581c752;
    ram_cell[     148] = 32'h0;  // 32'hace0830b;
    ram_cell[     149] = 32'h0;  // 32'hae53ca24;
    ram_cell[     150] = 32'h0;  // 32'hffb4b9cc;
    ram_cell[     151] = 32'h0;  // 32'h724bafcc;
    ram_cell[     152] = 32'h0;  // 32'h365acc78;
    ram_cell[     153] = 32'h0;  // 32'hdfac609e;
    ram_cell[     154] = 32'h0;  // 32'hdb1c3287;
    ram_cell[     155] = 32'h0;  // 32'h4d31ba88;
    ram_cell[     156] = 32'h0;  // 32'h25707ba6;
    ram_cell[     157] = 32'h0;  // 32'h8b3609f0;
    ram_cell[     158] = 32'h0;  // 32'hf6cb4815;
    ram_cell[     159] = 32'h0;  // 32'h4c8a829f;
    ram_cell[     160] = 32'h0;  // 32'h74b19b13;
    ram_cell[     161] = 32'h0;  // 32'h96bed440;
    ram_cell[     162] = 32'h0;  // 32'hdd1e78c9;
    ram_cell[     163] = 32'h0;  // 32'h0ba99ed5;
    ram_cell[     164] = 32'h0;  // 32'he8d9c5d5;
    ram_cell[     165] = 32'h0;  // 32'h41d5f3fd;
    ram_cell[     166] = 32'h0;  // 32'h7ff5dcff;
    ram_cell[     167] = 32'h0;  // 32'hd8db3019;
    ram_cell[     168] = 32'h0;  // 32'h26dbca89;
    ram_cell[     169] = 32'h0;  // 32'hbba55f4a;
    ram_cell[     170] = 32'h0;  // 32'hb6c32244;
    ram_cell[     171] = 32'h0;  // 32'hd8da35a0;
    ram_cell[     172] = 32'h0;  // 32'hcbdca60c;
    ram_cell[     173] = 32'h0;  // 32'hd9d02a25;
    ram_cell[     174] = 32'h0;  // 32'hbe3c3448;
    ram_cell[     175] = 32'h0;  // 32'he612a2b7;
    ram_cell[     176] = 32'h0;  // 32'h7cfef322;
    ram_cell[     177] = 32'h0;  // 32'hec3a5196;
    ram_cell[     178] = 32'h0;  // 32'h0fe9be65;
    ram_cell[     179] = 32'h0;  // 32'h78a16ef4;
    ram_cell[     180] = 32'h0;  // 32'h80a956e5;
    ram_cell[     181] = 32'h0;  // 32'h5d87e717;
    ram_cell[     182] = 32'h0;  // 32'h1e526cb5;
    ram_cell[     183] = 32'h0;  // 32'hc20d0ca1;
    ram_cell[     184] = 32'h0;  // 32'he933389b;
    ram_cell[     185] = 32'h0;  // 32'h79714e60;
    ram_cell[     186] = 32'h0;  // 32'h1f96f022;
    ram_cell[     187] = 32'h0;  // 32'h17a9fff0;
    ram_cell[     188] = 32'h0;  // 32'hab7b67c5;
    ram_cell[     189] = 32'h0;  // 32'h1896098b;
    ram_cell[     190] = 32'h0;  // 32'haf4b209a;
    ram_cell[     191] = 32'h0;  // 32'h0a6c7951;
    ram_cell[     192] = 32'h0;  // 32'hfd0a677c;
    ram_cell[     193] = 32'h0;  // 32'haf62012f;
    ram_cell[     194] = 32'h0;  // 32'hab287d02;
    ram_cell[     195] = 32'h0;  // 32'hf086e347;
    ram_cell[     196] = 32'h0;  // 32'h75c59aa7;
    ram_cell[     197] = 32'h0;  // 32'h57ef516a;
    ram_cell[     198] = 32'h0;  // 32'he890ace2;
    ram_cell[     199] = 32'h0;  // 32'h63e3dd59;
    ram_cell[     200] = 32'h0;  // 32'h707cc170;
    ram_cell[     201] = 32'h0;  // 32'h1d88912f;
    ram_cell[     202] = 32'h0;  // 32'h2c307ce2;
    ram_cell[     203] = 32'h0;  // 32'hd27c5397;
    ram_cell[     204] = 32'h0;  // 32'h48bec656;
    ram_cell[     205] = 32'h0;  // 32'h6386e30c;
    ram_cell[     206] = 32'h0;  // 32'h4425cc94;
    ram_cell[     207] = 32'h0;  // 32'he45d369d;
    ram_cell[     208] = 32'h0;  // 32'h95d5b13f;
    ram_cell[     209] = 32'h0;  // 32'h3ad6e27c;
    ram_cell[     210] = 32'h0;  // 32'h9c25013d;
    ram_cell[     211] = 32'h0;  // 32'h62899f7d;
    ram_cell[     212] = 32'h0;  // 32'he697f236;
    ram_cell[     213] = 32'h0;  // 32'h808d0bb1;
    ram_cell[     214] = 32'h0;  // 32'h599c2f3b;
    ram_cell[     215] = 32'h0;  // 32'h70f10031;
    ram_cell[     216] = 32'h0;  // 32'h7609abfc;
    ram_cell[     217] = 32'h0;  // 32'h571c30c5;
    ram_cell[     218] = 32'h0;  // 32'h611d8609;
    ram_cell[     219] = 32'h0;  // 32'h6f0a5699;
    ram_cell[     220] = 32'h0;  // 32'h02f954b0;
    ram_cell[     221] = 32'h0;  // 32'ha30247ae;
    ram_cell[     222] = 32'h0;  // 32'hb3032695;
    ram_cell[     223] = 32'h0;  // 32'h16c673bf;
    ram_cell[     224] = 32'h0;  // 32'h6300bbf8;
    ram_cell[     225] = 32'h0;  // 32'h66cace2b;
    ram_cell[     226] = 32'h0;  // 32'h3d8e2a75;
    ram_cell[     227] = 32'h0;  // 32'h66ba9362;
    ram_cell[     228] = 32'h0;  // 32'hb8464138;
    ram_cell[     229] = 32'h0;  // 32'hea5952e4;
    ram_cell[     230] = 32'h0;  // 32'hb019b9dd;
    ram_cell[     231] = 32'h0;  // 32'h35c93c5d;
    ram_cell[     232] = 32'h0;  // 32'ha2aefdac;
    ram_cell[     233] = 32'h0;  // 32'he98c34d1;
    ram_cell[     234] = 32'h0;  // 32'hec3087a3;
    ram_cell[     235] = 32'h0;  // 32'h6641b173;
    ram_cell[     236] = 32'h0;  // 32'hd9c28d85;
    ram_cell[     237] = 32'h0;  // 32'hf9a532db;
    ram_cell[     238] = 32'h0;  // 32'hea5b0dda;
    ram_cell[     239] = 32'h0;  // 32'hb863b59e;
    ram_cell[     240] = 32'h0;  // 32'h0442c678;
    ram_cell[     241] = 32'h0;  // 32'h3fd9b6b2;
    ram_cell[     242] = 32'h0;  // 32'ha0547bb4;
    ram_cell[     243] = 32'h0;  // 32'hffd7060d;
    ram_cell[     244] = 32'h0;  // 32'h534507a1;
    ram_cell[     245] = 32'h0;  // 32'h25d0ff5b;
    ram_cell[     246] = 32'h0;  // 32'hf79cb27a;
    ram_cell[     247] = 32'h0;  // 32'h2cb36cd1;
    ram_cell[     248] = 32'h0;  // 32'h8b6d9ad2;
    ram_cell[     249] = 32'h0;  // 32'h2f7fd078;
    ram_cell[     250] = 32'h0;  // 32'h648680cf;
    ram_cell[     251] = 32'h0;  // 32'hcb838cb4;
    ram_cell[     252] = 32'h0;  // 32'hb8c01765;
    ram_cell[     253] = 32'h0;  // 32'hc2a95efb;
    ram_cell[     254] = 32'h0;  // 32'ha11e31ed;
    ram_cell[     255] = 32'h0;  // 32'hb46c97f2;
    // src matrix A
    ram_cell[     256] = 32'h4fcea9ee;
    ram_cell[     257] = 32'ha3a0e92f;
    ram_cell[     258] = 32'ha9d3288e;
    ram_cell[     259] = 32'hd9b51570;
    ram_cell[     260] = 32'h8c85e200;
    ram_cell[     261] = 32'h2868d679;
    ram_cell[     262] = 32'h437c095f;
    ram_cell[     263] = 32'h7b8cbbca;
    ram_cell[     264] = 32'h45bf1abe;
    ram_cell[     265] = 32'ha2e7543b;
    ram_cell[     266] = 32'h99173ff3;
    ram_cell[     267] = 32'h20922af4;
    ram_cell[     268] = 32'h43341d0f;
    ram_cell[     269] = 32'hd04cb5e3;
    ram_cell[     270] = 32'h28f5a488;
    ram_cell[     271] = 32'h56f864b1;
    ram_cell[     272] = 32'h34f88154;
    ram_cell[     273] = 32'hb82a5465;
    ram_cell[     274] = 32'hf8acd4d9;
    ram_cell[     275] = 32'he7c54fe2;
    ram_cell[     276] = 32'h4e663589;
    ram_cell[     277] = 32'h6b158b21;
    ram_cell[     278] = 32'ha3b8a181;
    ram_cell[     279] = 32'h3fdd90d3;
    ram_cell[     280] = 32'h3b1aa920;
    ram_cell[     281] = 32'hcfe8fa3a;
    ram_cell[     282] = 32'h2990c54d;
    ram_cell[     283] = 32'hd17ef21c;
    ram_cell[     284] = 32'hb1287adb;
    ram_cell[     285] = 32'h35eb4963;
    ram_cell[     286] = 32'h2851d630;
    ram_cell[     287] = 32'h12afed26;
    ram_cell[     288] = 32'h7e375d7b;
    ram_cell[     289] = 32'h1322ff81;
    ram_cell[     290] = 32'h65ee81b3;
    ram_cell[     291] = 32'hcbe674aa;
    ram_cell[     292] = 32'h775c6bb0;
    ram_cell[     293] = 32'h260c1794;
    ram_cell[     294] = 32'h9f87375d;
    ram_cell[     295] = 32'h3ee89055;
    ram_cell[     296] = 32'h09bd85a0;
    ram_cell[     297] = 32'he6f05e9a;
    ram_cell[     298] = 32'h753270b8;
    ram_cell[     299] = 32'h71bb991f;
    ram_cell[     300] = 32'hf3177fd2;
    ram_cell[     301] = 32'hb0dc9868;
    ram_cell[     302] = 32'h5aa7750b;
    ram_cell[     303] = 32'he1662657;
    ram_cell[     304] = 32'h61e2162d;
    ram_cell[     305] = 32'hbc166a6d;
    ram_cell[     306] = 32'h088eea5d;
    ram_cell[     307] = 32'h21e9be72;
    ram_cell[     308] = 32'hd37ea0b2;
    ram_cell[     309] = 32'h8b58ea9f;
    ram_cell[     310] = 32'h4c5425bc;
    ram_cell[     311] = 32'h64202c18;
    ram_cell[     312] = 32'hcc8ee3ca;
    ram_cell[     313] = 32'h7d3aff5d;
    ram_cell[     314] = 32'hc1a31542;
    ram_cell[     315] = 32'hd980d20b;
    ram_cell[     316] = 32'h1697e038;
    ram_cell[     317] = 32'haf64bb96;
    ram_cell[     318] = 32'h87dda48c;
    ram_cell[     319] = 32'h34a7f355;
    ram_cell[     320] = 32'h10c2cc2a;
    ram_cell[     321] = 32'h4de87d07;
    ram_cell[     322] = 32'he06127ce;
    ram_cell[     323] = 32'h15b07c03;
    ram_cell[     324] = 32'h5161dfc6;
    ram_cell[     325] = 32'ha1f2f5bf;
    ram_cell[     326] = 32'ha165c6fd;
    ram_cell[     327] = 32'hdfe58f70;
    ram_cell[     328] = 32'h6fec28b9;
    ram_cell[     329] = 32'h71d582f4;
    ram_cell[     330] = 32'h81a347d9;
    ram_cell[     331] = 32'h4166d94b;
    ram_cell[     332] = 32'he56c5190;
    ram_cell[     333] = 32'he9c0a42a;
    ram_cell[     334] = 32'hb65383d9;
    ram_cell[     335] = 32'hd7096005;
    ram_cell[     336] = 32'h66634f3c;
    ram_cell[     337] = 32'h16f26fd1;
    ram_cell[     338] = 32'hb5ca0b67;
    ram_cell[     339] = 32'he0d29882;
    ram_cell[     340] = 32'hb6cb9867;
    ram_cell[     341] = 32'h6d1dd730;
    ram_cell[     342] = 32'h88eb71d4;
    ram_cell[     343] = 32'h13a698d5;
    ram_cell[     344] = 32'h9d5c893b;
    ram_cell[     345] = 32'h2e7e70ec;
    ram_cell[     346] = 32'h6d925d49;
    ram_cell[     347] = 32'h7098945f;
    ram_cell[     348] = 32'hdf301a5e;
    ram_cell[     349] = 32'hb76cc515;
    ram_cell[     350] = 32'h917129ed;
    ram_cell[     351] = 32'h89adabb7;
    ram_cell[     352] = 32'h73594c32;
    ram_cell[     353] = 32'h8507c7a0;
    ram_cell[     354] = 32'hea3d663c;
    ram_cell[     355] = 32'hd684a414;
    ram_cell[     356] = 32'h62f8c211;
    ram_cell[     357] = 32'h82adab0c;
    ram_cell[     358] = 32'hb714fcc9;
    ram_cell[     359] = 32'hf0882e8f;
    ram_cell[     360] = 32'h6dd7aa54;
    ram_cell[     361] = 32'h5552303a;
    ram_cell[     362] = 32'h2948884f;
    ram_cell[     363] = 32'h93ce78b0;
    ram_cell[     364] = 32'h6ab10b1e;
    ram_cell[     365] = 32'h7c13a53a;
    ram_cell[     366] = 32'h25bd8526;
    ram_cell[     367] = 32'h4f8dd5c7;
    ram_cell[     368] = 32'hd6e892df;
    ram_cell[     369] = 32'h90787009;
    ram_cell[     370] = 32'h1453aea9;
    ram_cell[     371] = 32'h602955cf;
    ram_cell[     372] = 32'hd3a98d63;
    ram_cell[     373] = 32'hf130b6aa;
    ram_cell[     374] = 32'h79afc01e;
    ram_cell[     375] = 32'h1234b49b;
    ram_cell[     376] = 32'hf3fe6083;
    ram_cell[     377] = 32'hd7b00602;
    ram_cell[     378] = 32'h681c106a;
    ram_cell[     379] = 32'hc8049906;
    ram_cell[     380] = 32'h40d36274;
    ram_cell[     381] = 32'hc2581ac4;
    ram_cell[     382] = 32'h2b2b5eb3;
    ram_cell[     383] = 32'hfa2f673b;
    ram_cell[     384] = 32'hac022359;
    ram_cell[     385] = 32'h97f4d5f4;
    ram_cell[     386] = 32'hb124da56;
    ram_cell[     387] = 32'h01f3d711;
    ram_cell[     388] = 32'h040a7995;
    ram_cell[     389] = 32'h8ceddf45;
    ram_cell[     390] = 32'hdc70f18b;
    ram_cell[     391] = 32'h6be9eb7f;
    ram_cell[     392] = 32'h7978baeb;
    ram_cell[     393] = 32'h70e883df;
    ram_cell[     394] = 32'hae467252;
    ram_cell[     395] = 32'hf95e2186;
    ram_cell[     396] = 32'h542d88a2;
    ram_cell[     397] = 32'h575ec93e;
    ram_cell[     398] = 32'h66475c60;
    ram_cell[     399] = 32'h64db5f4a;
    ram_cell[     400] = 32'hc1ea12b0;
    ram_cell[     401] = 32'h5c26f2be;
    ram_cell[     402] = 32'h85326f0b;
    ram_cell[     403] = 32'h5f7a5168;
    ram_cell[     404] = 32'h771b62bf;
    ram_cell[     405] = 32'hf06a504a;
    ram_cell[     406] = 32'h16196ccb;
    ram_cell[     407] = 32'hf8e40081;
    ram_cell[     408] = 32'hcf486a84;
    ram_cell[     409] = 32'hc9e85394;
    ram_cell[     410] = 32'h92462d5d;
    ram_cell[     411] = 32'hacaf8b3a;
    ram_cell[     412] = 32'habbeceed;
    ram_cell[     413] = 32'h73917ea8;
    ram_cell[     414] = 32'h92ad0bb2;
    ram_cell[     415] = 32'h7ab10d4e;
    ram_cell[     416] = 32'h906e31d4;
    ram_cell[     417] = 32'hbb12cc5f;
    ram_cell[     418] = 32'h19794564;
    ram_cell[     419] = 32'ha010e87e;
    ram_cell[     420] = 32'heb072e3a;
    ram_cell[     421] = 32'h453b11f2;
    ram_cell[     422] = 32'hc218d31c;
    ram_cell[     423] = 32'hba06cb49;
    ram_cell[     424] = 32'hec93c67f;
    ram_cell[     425] = 32'hbe5f0086;
    ram_cell[     426] = 32'h905abebe;
    ram_cell[     427] = 32'hfb3bc3ad;
    ram_cell[     428] = 32'h3ce8fd92;
    ram_cell[     429] = 32'h303decfd;
    ram_cell[     430] = 32'h25c4447b;
    ram_cell[     431] = 32'hfd5487d6;
    ram_cell[     432] = 32'hc824316a;
    ram_cell[     433] = 32'h4dbaebd4;
    ram_cell[     434] = 32'h1341d3de;
    ram_cell[     435] = 32'h18ea62cf;
    ram_cell[     436] = 32'hc09ac163;
    ram_cell[     437] = 32'h2458831d;
    ram_cell[     438] = 32'hf8cf1238;
    ram_cell[     439] = 32'haf514cf9;
    ram_cell[     440] = 32'hb8568908;
    ram_cell[     441] = 32'h653429c2;
    ram_cell[     442] = 32'ha93cba02;
    ram_cell[     443] = 32'hae5b5106;
    ram_cell[     444] = 32'hc780647a;
    ram_cell[     445] = 32'hd77dd152;
    ram_cell[     446] = 32'h2919525c;
    ram_cell[     447] = 32'h43b154b6;
    ram_cell[     448] = 32'h1b91edd3;
    ram_cell[     449] = 32'hfe36e52c;
    ram_cell[     450] = 32'h52350c61;
    ram_cell[     451] = 32'h9660b47e;
    ram_cell[     452] = 32'h258b4db1;
    ram_cell[     453] = 32'hddc43bfa;
    ram_cell[     454] = 32'h4acaf3c1;
    ram_cell[     455] = 32'hb63f756b;
    ram_cell[     456] = 32'h63c53e91;
    ram_cell[     457] = 32'h8ab3f9b7;
    ram_cell[     458] = 32'h72a03235;
    ram_cell[     459] = 32'h9e2fac96;
    ram_cell[     460] = 32'he72f098c;
    ram_cell[     461] = 32'h4a219948;
    ram_cell[     462] = 32'h9f72c9ee;
    ram_cell[     463] = 32'hae766f9a;
    ram_cell[     464] = 32'h884846f6;
    ram_cell[     465] = 32'hdaa042e1;
    ram_cell[     466] = 32'hb22b03b4;
    ram_cell[     467] = 32'h61f9cce3;
    ram_cell[     468] = 32'hf9795d9d;
    ram_cell[     469] = 32'h5922defe;
    ram_cell[     470] = 32'h9ddf961c;
    ram_cell[     471] = 32'h5bd0eafc;
    ram_cell[     472] = 32'h4ad796e4;
    ram_cell[     473] = 32'he69723d2;
    ram_cell[     474] = 32'ha3c6b333;
    ram_cell[     475] = 32'h64e0010c;
    ram_cell[     476] = 32'hde284f0c;
    ram_cell[     477] = 32'hff9dbb5f;
    ram_cell[     478] = 32'h4aaf5aed;
    ram_cell[     479] = 32'h8d578bf2;
    ram_cell[     480] = 32'h8f11cdea;
    ram_cell[     481] = 32'he307bd0f;
    ram_cell[     482] = 32'h42615389;
    ram_cell[     483] = 32'h083cf57e;
    ram_cell[     484] = 32'h363cee77;
    ram_cell[     485] = 32'he719cc6c;
    ram_cell[     486] = 32'h5e79ce20;
    ram_cell[     487] = 32'h3c8ce626;
    ram_cell[     488] = 32'h63e0346e;
    ram_cell[     489] = 32'h1c251c7d;
    ram_cell[     490] = 32'h825d2f6c;
    ram_cell[     491] = 32'hf25a435d;
    ram_cell[     492] = 32'h8db6264f;
    ram_cell[     493] = 32'h9d294545;
    ram_cell[     494] = 32'hfe746f85;
    ram_cell[     495] = 32'h2a0142be;
    ram_cell[     496] = 32'h06050025;
    ram_cell[     497] = 32'h82282628;
    ram_cell[     498] = 32'h911478d3;
    ram_cell[     499] = 32'hcf8f43e9;
    ram_cell[     500] = 32'hb2863968;
    ram_cell[     501] = 32'h601d3324;
    ram_cell[     502] = 32'haab0911b;
    ram_cell[     503] = 32'hc2c82030;
    ram_cell[     504] = 32'h343b0f81;
    ram_cell[     505] = 32'h24c14e85;
    ram_cell[     506] = 32'h0d6698fc;
    ram_cell[     507] = 32'hd3762955;
    ram_cell[     508] = 32'hd2c5fbe5;
    ram_cell[     509] = 32'h5d694a5b;
    ram_cell[     510] = 32'h2bc463b5;
    ram_cell[     511] = 32'he78e4525;
    // src matrix B
    ram_cell[     512] = 32'hccf62842;
    ram_cell[     513] = 32'h101ca672;
    ram_cell[     514] = 32'h3a0e4eb9;
    ram_cell[     515] = 32'h5cefacf4;
    ram_cell[     516] = 32'hd594d9ad;
    ram_cell[     517] = 32'h46d558f8;
    ram_cell[     518] = 32'h1ae6bf5f;
    ram_cell[     519] = 32'h7236426c;
    ram_cell[     520] = 32'h5ba3d872;
    ram_cell[     521] = 32'h236f0dd3;
    ram_cell[     522] = 32'hfc9cb741;
    ram_cell[     523] = 32'h9903468e;
    ram_cell[     524] = 32'h6da6399a;
    ram_cell[     525] = 32'h338df8ea;
    ram_cell[     526] = 32'h27881512;
    ram_cell[     527] = 32'hcaf1bfcd;
    ram_cell[     528] = 32'hecf8299c;
    ram_cell[     529] = 32'hd79e3119;
    ram_cell[     530] = 32'h3f7bc7f0;
    ram_cell[     531] = 32'h6718c902;
    ram_cell[     532] = 32'hf68d49d6;
    ram_cell[     533] = 32'h856b957f;
    ram_cell[     534] = 32'h1ac2646b;
    ram_cell[     535] = 32'h4e979faf;
    ram_cell[     536] = 32'hf72587c2;
    ram_cell[     537] = 32'h4ad903d7;
    ram_cell[     538] = 32'h81cedb03;
    ram_cell[     539] = 32'h38d44f31;
    ram_cell[     540] = 32'h3f27928a;
    ram_cell[     541] = 32'h2c05fa67;
    ram_cell[     542] = 32'h45436f11;
    ram_cell[     543] = 32'h6609c0f6;
    ram_cell[     544] = 32'h85ffdf43;
    ram_cell[     545] = 32'hbe014154;
    ram_cell[     546] = 32'he71e87fc;
    ram_cell[     547] = 32'h660bd0e4;
    ram_cell[     548] = 32'hd09d6aca;
    ram_cell[     549] = 32'h38e23737;
    ram_cell[     550] = 32'h82579ce0;
    ram_cell[     551] = 32'hf2e5cfef;
    ram_cell[     552] = 32'h9a982ba8;
    ram_cell[     553] = 32'hc009f126;
    ram_cell[     554] = 32'h78a79b6c;
    ram_cell[     555] = 32'haa7de6f4;
    ram_cell[     556] = 32'hb5675589;
    ram_cell[     557] = 32'h4a523e77;
    ram_cell[     558] = 32'h4d3bb499;
    ram_cell[     559] = 32'hc3bf301b;
    ram_cell[     560] = 32'hadc17307;
    ram_cell[     561] = 32'h027a7f79;
    ram_cell[     562] = 32'hffd3ae70;
    ram_cell[     563] = 32'h2aef16f5;
    ram_cell[     564] = 32'h647019da;
    ram_cell[     565] = 32'h6aae27ba;
    ram_cell[     566] = 32'h38e2acb8;
    ram_cell[     567] = 32'h46636ce2;
    ram_cell[     568] = 32'h286bd65a;
    ram_cell[     569] = 32'h9e9c4e98;
    ram_cell[     570] = 32'h0f975f0d;
    ram_cell[     571] = 32'h50ce6072;
    ram_cell[     572] = 32'h33acf38f;
    ram_cell[     573] = 32'hbf214ee7;
    ram_cell[     574] = 32'h314b9771;
    ram_cell[     575] = 32'h6046abba;
    ram_cell[     576] = 32'hef13928e;
    ram_cell[     577] = 32'h098ed21a;
    ram_cell[     578] = 32'h526b1816;
    ram_cell[     579] = 32'h29d20365;
    ram_cell[     580] = 32'h0a2fe9c2;
    ram_cell[     581] = 32'h1e36f76b;
    ram_cell[     582] = 32'h9d11b3f8;
    ram_cell[     583] = 32'he948c1ab;
    ram_cell[     584] = 32'h6e18f540;
    ram_cell[     585] = 32'hf32833ee;
    ram_cell[     586] = 32'h7134bd23;
    ram_cell[     587] = 32'hbd12ce9d;
    ram_cell[     588] = 32'h80af3bb5;
    ram_cell[     589] = 32'h30bfb85d;
    ram_cell[     590] = 32'h245dded4;
    ram_cell[     591] = 32'h6d76f608;
    ram_cell[     592] = 32'h65c20153;
    ram_cell[     593] = 32'h622c4dcb;
    ram_cell[     594] = 32'hdd0d8401;
    ram_cell[     595] = 32'h5ab1520b;
    ram_cell[     596] = 32'hc17cb9bf;
    ram_cell[     597] = 32'h8aa8f26f;
    ram_cell[     598] = 32'ha6532c2e;
    ram_cell[     599] = 32'h0b9a13b3;
    ram_cell[     600] = 32'hd0e34cda;
    ram_cell[     601] = 32'h027cd757;
    ram_cell[     602] = 32'hf5d0fde8;
    ram_cell[     603] = 32'h3c22cbb6;
    ram_cell[     604] = 32'h18a88cf4;
    ram_cell[     605] = 32'h1ce9afe5;
    ram_cell[     606] = 32'h9bc36e49;
    ram_cell[     607] = 32'h4f697e50;
    ram_cell[     608] = 32'hdb4703ce;
    ram_cell[     609] = 32'hd6d77063;
    ram_cell[     610] = 32'hc021f1c4;
    ram_cell[     611] = 32'hf7874cf3;
    ram_cell[     612] = 32'h4e17315d;
    ram_cell[     613] = 32'h2dc8f7ce;
    ram_cell[     614] = 32'h29b741e2;
    ram_cell[     615] = 32'h31c12ccf;
    ram_cell[     616] = 32'h82f7cf56;
    ram_cell[     617] = 32'hf50e8642;
    ram_cell[     618] = 32'h6d5d4302;
    ram_cell[     619] = 32'h92d63e36;
    ram_cell[     620] = 32'h0915cc27;
    ram_cell[     621] = 32'h0349a677;
    ram_cell[     622] = 32'h89bbd4fd;
    ram_cell[     623] = 32'h28fda011;
    ram_cell[     624] = 32'h8920f2ce;
    ram_cell[     625] = 32'hc6c0f492;
    ram_cell[     626] = 32'h5ba6bf5a;
    ram_cell[     627] = 32'h58e0b725;
    ram_cell[     628] = 32'h8376b868;
    ram_cell[     629] = 32'h5e61ba49;
    ram_cell[     630] = 32'hf4ef6b57;
    ram_cell[     631] = 32'h0b5dc851;
    ram_cell[     632] = 32'h645dfbd1;
    ram_cell[     633] = 32'h4e7b2c9f;
    ram_cell[     634] = 32'hc7ed7702;
    ram_cell[     635] = 32'h47c89eaf;
    ram_cell[     636] = 32'h8b0a4575;
    ram_cell[     637] = 32'ha289ce44;
    ram_cell[     638] = 32'hb8d76c5e;
    ram_cell[     639] = 32'h5dc965db;
    ram_cell[     640] = 32'h07078b2f;
    ram_cell[     641] = 32'h5c8e60a7;
    ram_cell[     642] = 32'hb398a2c2;
    ram_cell[     643] = 32'he658e2cf;
    ram_cell[     644] = 32'h0f8ec3c5;
    ram_cell[     645] = 32'hb634ea7b;
    ram_cell[     646] = 32'h6e84c2af;
    ram_cell[     647] = 32'h8febcd27;
    ram_cell[     648] = 32'he85627d8;
    ram_cell[     649] = 32'h799fa5fb;
    ram_cell[     650] = 32'h57dbf399;
    ram_cell[     651] = 32'h0b01ad3b;
    ram_cell[     652] = 32'ha72e43ac;
    ram_cell[     653] = 32'h5b6ea1de;
    ram_cell[     654] = 32'hdcf6d04f;
    ram_cell[     655] = 32'h6d67a45b;
    ram_cell[     656] = 32'h23a0de9c;
    ram_cell[     657] = 32'h4b8e4d79;
    ram_cell[     658] = 32'h9e343e84;
    ram_cell[     659] = 32'hd437e6a8;
    ram_cell[     660] = 32'hf01c3336;
    ram_cell[     661] = 32'h0a073b58;
    ram_cell[     662] = 32'h408c20c4;
    ram_cell[     663] = 32'h6a348a5e;
    ram_cell[     664] = 32'hc1cab22d;
    ram_cell[     665] = 32'h5e04a3a8;
    ram_cell[     666] = 32'h1073d3ad;
    ram_cell[     667] = 32'h216e78f6;
    ram_cell[     668] = 32'h376c2945;
    ram_cell[     669] = 32'hbfe68203;
    ram_cell[     670] = 32'hc2f68c47;
    ram_cell[     671] = 32'hf567250c;
    ram_cell[     672] = 32'h5e999c4c;
    ram_cell[     673] = 32'h3cb9e69c;
    ram_cell[     674] = 32'h951b9861;
    ram_cell[     675] = 32'h98915991;
    ram_cell[     676] = 32'hae07b314;
    ram_cell[     677] = 32'h299f2888;
    ram_cell[     678] = 32'h9f733bc3;
    ram_cell[     679] = 32'h1c9507d0;
    ram_cell[     680] = 32'h6d9f5e32;
    ram_cell[     681] = 32'h55fb1f04;
    ram_cell[     682] = 32'hfdfb0cf6;
    ram_cell[     683] = 32'haa4a6228;
    ram_cell[     684] = 32'h8264ec55;
    ram_cell[     685] = 32'h39eca3dc;
    ram_cell[     686] = 32'h4101d1e0;
    ram_cell[     687] = 32'h925ab926;
    ram_cell[     688] = 32'h5865ef10;
    ram_cell[     689] = 32'h1525e71e;
    ram_cell[     690] = 32'h47d81447;
    ram_cell[     691] = 32'hbcad219b;
    ram_cell[     692] = 32'h4bb2e5b6;
    ram_cell[     693] = 32'hb36d53d3;
    ram_cell[     694] = 32'hb49136b7;
    ram_cell[     695] = 32'h1206efa3;
    ram_cell[     696] = 32'he89bd1d2;
    ram_cell[     697] = 32'hd9f359b5;
    ram_cell[     698] = 32'h4a12e2ca;
    ram_cell[     699] = 32'h4d7b09b0;
    ram_cell[     700] = 32'h2c85c574;
    ram_cell[     701] = 32'h7869c69d;
    ram_cell[     702] = 32'h3e1d95df;
    ram_cell[     703] = 32'h2a797d9c;
    ram_cell[     704] = 32'h05eff791;
    ram_cell[     705] = 32'hba855dc5;
    ram_cell[     706] = 32'h406b97c4;
    ram_cell[     707] = 32'h6f1d72e4;
    ram_cell[     708] = 32'h339bcfb8;
    ram_cell[     709] = 32'h0c730c63;
    ram_cell[     710] = 32'he1d80758;
    ram_cell[     711] = 32'hbde4e434;
    ram_cell[     712] = 32'hf80aef71;
    ram_cell[     713] = 32'h97ca8eff;
    ram_cell[     714] = 32'hda42fe32;
    ram_cell[     715] = 32'h1fa245f2;
    ram_cell[     716] = 32'h336ce2af;
    ram_cell[     717] = 32'hb5bf1241;
    ram_cell[     718] = 32'ha13aa579;
    ram_cell[     719] = 32'h56c952d8;
    ram_cell[     720] = 32'hd6ce7918;
    ram_cell[     721] = 32'hfbc2b69e;
    ram_cell[     722] = 32'h1afd7d12;
    ram_cell[     723] = 32'h67b21c39;
    ram_cell[     724] = 32'h16374bc7;
    ram_cell[     725] = 32'h0d362b83;
    ram_cell[     726] = 32'he084d279;
    ram_cell[     727] = 32'h8cc1e045;
    ram_cell[     728] = 32'hff8a3925;
    ram_cell[     729] = 32'h820d72db;
    ram_cell[     730] = 32'h48bf99e4;
    ram_cell[     731] = 32'h50dc22c0;
    ram_cell[     732] = 32'h6ac1886c;
    ram_cell[     733] = 32'h1511fe91;
    ram_cell[     734] = 32'h7c917cc4;
    ram_cell[     735] = 32'he1f31247;
    ram_cell[     736] = 32'h099d5dca;
    ram_cell[     737] = 32'h42f2df80;
    ram_cell[     738] = 32'h55433ebe;
    ram_cell[     739] = 32'h04344d55;
    ram_cell[     740] = 32'he9dd0be5;
    ram_cell[     741] = 32'h82dcd2cc;
    ram_cell[     742] = 32'hed60dcfc;
    ram_cell[     743] = 32'h3a807f60;
    ram_cell[     744] = 32'h19e5cc41;
    ram_cell[     745] = 32'h4de8c557;
    ram_cell[     746] = 32'h614baaee;
    ram_cell[     747] = 32'h46743e65;
    ram_cell[     748] = 32'haf318fa9;
    ram_cell[     749] = 32'ha2d41c2a;
    ram_cell[     750] = 32'h4983e89f;
    ram_cell[     751] = 32'h521ddacc;
    ram_cell[     752] = 32'h8e24e930;
    ram_cell[     753] = 32'h6dcd467d;
    ram_cell[     754] = 32'h68ad810a;
    ram_cell[     755] = 32'h64714203;
    ram_cell[     756] = 32'h7f096bb8;
    ram_cell[     757] = 32'hf7c66a40;
    ram_cell[     758] = 32'he5965a7a;
    ram_cell[     759] = 32'h863ca4ec;
    ram_cell[     760] = 32'h258091f2;
    ram_cell[     761] = 32'hf9380800;
    ram_cell[     762] = 32'hbec93c55;
    ram_cell[     763] = 32'hb6c4ad1a;
    ram_cell[     764] = 32'h5d1ceea1;
    ram_cell[     765] = 32'h3d8387ec;
    ram_cell[     766] = 32'h62151fbb;
    ram_cell[     767] = 32'h4cf429a5;
end

endmodule

