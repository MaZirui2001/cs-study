// asm file name: bht.S
module InstructionCache(
    input wire clk,
    input wire write_en,
    input wire [31:2] addr, debug_addr,
    input wire [31:0] debug_input,
    output reg [31:0] data, debug_data
);

    // local variable
    wire addr_valid = (addr[31:14] == 18'h0);
    wire debug_addr_valid = (debug_addr[31:14] == 18'h0);
    wire [11:0] dealt_addr = addr[13:2];
    wire [11:0] dealt_debug_addr = debug_addr[13:2];
    // cache content
    reg [31:0] inst_cache[0:4095];


    initial begin
        data = 32'h0;
        debug_data = 32'h0;
        inst_cache[       0] = 32'h00000293;
        inst_cache[       1] = 32'h00000313;
        inst_cache[       2] = 32'h00000393;
        inst_cache[       3] = 32'h00a00e13;
        inst_cache[       4] = 32'h00138393;
        inst_cache[       5] = 32'h00530333;
        inst_cache[       6] = 32'h00128293;
        inst_cache[       7] = 32'hffc29ce3;
        inst_cache[       8] = 32'h00000293;
        inst_cache[       9] = 32'hffc396e3;
        inst_cache[      10] = 32'h00130313;
        inst_cache[      11] = 32'h0000006f;
end

    always@(posedge clk)
    begin
        data <= addr_valid ? inst_cache[dealt_addr] : 32'h0;
        debug_data <= debug_addr_valid ? inst_cache[dealt_debug_addr] : 32'h0;
        if(write_en & debug_addr_valid) 
            inst_cache[dealt_debug_addr] <= debug_input;
    end

endmodule
